`timescale 1ns / 1ps

module SytemZ_3(

    );
endmodule
